`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/04/14 17:23:31
// Design Name: 
// Module Name: draw_board
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module draw_board(
    input [3:0]r, g, b,
    input [3:0]dirc,
    input draw,
    output [3:0]disr, disg, disb,
    output hs, vs
    );
endmodule
